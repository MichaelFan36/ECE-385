module testbench2();

timeunit 10ns;

timeprecision 1ns;

logic Clk;

logic [9:0] SW;

logic Run, Continue;

logic [9:0] LED;

logic [6:0] HEX0, HEX1, HEX2, HEX3;

logic [6:0] HEX0_, HEX1_, HEX2_, HEX3_;

integer ErrorCnt = 0;



slc3_testtop tp(.*);

//****     ***** **** *** ***  ***
//********   *****   ******    ***
//****   *****   ****    **   *  *     
//************   ********  *** ***
//*** *** **  *****   ***** ******
//*** ***** **  ***   ***** ** ***
//**  **  ** ** ***  *** ** *  ***
//*************   ****************
	

always begin : CLOCK_GENERATION
#1 Clk = ~Clk;
end

initial begin: CLOCK_INITIALIZATION
    Clk = 0;
end 

initial begin: TEST_VECTORS
Run = 1'b1; 
Continue = 1'b1;


// initialize test case
SW = 10'b0000000011;				// test 1
//SW = 10'b0000000110;				// test 2
//SW = 10'b0000001100;				// test 3
//SW = 10'b0000010100;				// test 4
//SW = 10'b0000110001;				// test 5
//SW = 10'b0000101010;					// test 6

// reset
#2 Run = 0;
#2 Continue = 0;
#20 Run = 1;
#20 Continue = 1;

#2 Run = 0;//triger Run
#2 Run = 1;

//// test 1
#100 SW = 10'b0000110011;

#100 SW = 10'b0100110011;

#100 SW = 10'b0101010101;
////

//// test 2
//#100 SW = 10'b0000110011;
//
//#10 Continue = 0;
//#20 Continue = 1;
//
//#100 SW = 10'b0100110011;
//
//#10 Continue = 0;
//#20 Continue = 1;
//
//#100 SW = 10'b0101010101;
//
//#10 Continue = 0;
//#20 Continue = 1;
////

//// test 3
//#300 Continue = 0;
//#20 Continue = 1;
//
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
////

//// test 4
//
//#300 SW = 10'b1011110010;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 SW = 10'b1101001010;
//
//#300 Continue = 0;
//#20 Continue = 1;
//// result should be SW = 10'b01 1011 1000;
//


// test 5

//#300 SW = 10'b0000000011; // 3
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 SW = 10'b0000000100; // 4
//
//#300 Continue = 0;
//#20 Continue = 1;
//// result should be SW = 10'b0000 0000 1100;
//
//#1000 ;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 SW = 10'b0000000011; // 3
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 SW = 10'b0000000101; // 5
//
//#300 Continue = 0;
//#20 Continue = 1;
// result should be SW = 10'b0000 0000 1111;

// test 7
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
//
//#300 Continue = 0;
//#20 Continue = 1;
end

endmodule
